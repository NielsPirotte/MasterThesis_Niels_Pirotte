p50 vhdl ref manual
